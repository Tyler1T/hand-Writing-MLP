module neuron(input bias[15:0] );
    for(int i = 0; i < )

endmodule // neuron

module network (data, result);
    input logic [0:15] data [783:0];
    output logic [0:15] result[9:0];
    wire [0:15] layer1_output[199:0];
    wire [0:15] layer2_output[49:0];

    neuron_layer1 n1_0 (data, 0, layer1_output[0]);
    neuron_layer1 n1_1 (data, 1, layer1_output[1]);
    neuron_layer1 n1_2 (data, 2, layer1_output[2]);
    neuron_layer1 n1_3 (data, 3, layer1_output[3]);
    neuron_layer1 n1_4 (data, 4, layer1_output[4]);
    neuron_layer1 n1_5 (data, 5, layer1_output[5]);
    neuron_layer1 n1_6 (data, 6, layer1_output[6]);
    neuron_layer1 n1_7 (data, 7, layer1_output[7]);
    neuron_layer1 n1_8 (data, 8, layer1_output[8]);
    neuron_layer1 n1_9 (data, 9, layer1_output[9]);
    neuron_layer1 n1_10 (data, 10, layer1_output[10]);
    neuron_layer1 n1_11 (data, 11, layer1_output[11]);
    neuron_layer1 n1_12 (data, 12, layer1_output[12]);
    neuron_layer1 n1_13 (data, 13, layer1_output[13]);
    neuron_layer1 n1_14 (data, 14, layer1_output[14]);
    neuron_layer1 n1_15 (data, 15, layer1_output[15]);
    neuron_layer1 n1_16 (data, 16, layer1_output[16]);
    neuron_layer1 n1_17 (data, 17, layer1_output[17]);
    neuron_layer1 n1_18 (data, 18, layer1_output[18]);
    neuron_layer1 n1_19 (data, 19, layer1_output[19]);
    neuron_layer1 n1_20 (data, 20, layer1_output[20]);
    neuron_layer1 n1_21 (data, 21, layer1_output[21]);
    neuron_layer1 n1_22 (data, 22, layer1_output[22]);
    neuron_layer1 n1_23 (data, 23, layer1_output[23]);
    neuron_layer1 n1_24 (data, 24, layer1_output[24]);
    neuron_layer1 n1_25 (data, 25, layer1_output[25]);
    neuron_layer1 n1_26 (data, 26, layer1_output[26]);
    neuron_layer1 n1_27 (data, 27, layer1_output[27]);
    neuron_layer1 n1_28 (data, 28, layer1_output[28]);
    neuron_layer1 n1_29 (data, 29, layer1_output[29]);
    neuron_layer1 n1_30 (data, 30, layer1_output[30]);
    neuron_layer1 n1_31 (data, 31, layer1_output[31]);
    neuron_layer1 n1_32 (data, 32, layer1_output[32]);
    neuron_layer1 n1_33 (data, 33, layer1_output[33]);
    neuron_layer1 n1_34 (data, 34, layer1_output[34]);
    neuron_layer1 n1_35 (data, 35, layer1_output[35]);
    neuron_layer1 n1_36 (data, 36, layer1_output[36]);
    neuron_layer1 n1_37 (data, 37, layer1_output[37]);
    neuron_layer1 n1_38 (data, 38, layer1_output[38]);
    neuron_layer1 n1_39 (data, 39, layer1_output[39]);
    neuron_layer1 n1_40 (data, 40, layer1_output[40]);
    neuron_layer1 n1_41 (data, 41, layer1_output[41]);
    neuron_layer1 n1_42 (data, 42, layer1_output[42]);
    neuron_layer1 n1_43 (data, 43, layer1_output[43]);
    neuron_layer1 n1_44 (data, 44, layer1_output[44]);
    neuron_layer1 n1_45 (data, 45, layer1_output[45]);
    neuron_layer1 n1_46 (data, 46, layer1_output[46]);
    neuron_layer1 n1_47 (data, 47, layer1_output[47]);
    neuron_layer1 n1_48 (data, 48, layer1_output[48]);
    neuron_layer1 n1_49 (data, 49, layer1_output[49]);
    neuron_layer1 n1_50 (data, 50, layer1_output[50]);
    neuron_layer1 n1_51 (data, 51, layer1_output[51]);
    neuron_layer1 n1_52 (data, 52, layer1_output[52]);
    neuron_layer1 n1_53 (data, 53, layer1_output[53]);
    neuron_layer1 n1_54 (data, 54, layer1_output[54]);
    neuron_layer1 n1_55 (data, 55, layer1_output[55]);
    neuron_layer1 n1_56 (data, 56, layer1_output[56]);
    neuron_layer1 n1_57 (data, 57, layer1_output[57]);
    neuron_layer1 n1_58 (data, 58, layer1_output[58]);
    neuron_layer1 n1_59 (data, 59, layer1_output[59]);
    neuron_layer1 n1_60 (data, 60, layer1_output[60]);
    neuron_layer1 n1_61 (data, 61, layer1_output[61]);
    neuron_layer1 n1_62 (data, 62, layer1_output[62]);
    neuron_layer1 n1_63 (data, 63, layer1_output[63]);
    neuron_layer1 n1_64 (data, 64, layer1_output[64]);
    neuron_layer1 n1_65 (data, 65, layer1_output[65]);
    neuron_layer1 n1_66 (data, 66, layer1_output[66]);
    neuron_layer1 n1_67 (data, 67, layer1_output[67]);
    neuron_layer1 n1_68 (data, 68, layer1_output[68]);
    neuron_layer1 n1_69 (data, 69, layer1_output[69]);
    neuron_layer1 n1_70 (data, 70, layer1_output[70]);
    neuron_layer1 n1_71 (data, 71, layer1_output[71]);
    neuron_layer1 n1_72 (data, 72, layer1_output[72]);
    neuron_layer1 n1_73 (data, 73, layer1_output[73]);
    neuron_layer1 n1_74 (data, 74, layer1_output[74]);
    neuron_layer1 n1_75 (data, 75, layer1_output[75]);
    neuron_layer1 n1_76 (data, 76, layer1_output[76]);
    neuron_layer1 n1_77 (data, 77, layer1_output[77]);
    neuron_layer1 n1_78 (data, 78, layer1_output[78]);
    neuron_layer1 n1_79 (data, 79, layer1_output[79]);
    neuron_layer1 n1_80 (data, 80, layer1_output[80]);
    neuron_layer1 n1_81 (data, 81, layer1_output[81]);
    neuron_layer1 n1_82 (data, 82, layer1_output[82]);
    neuron_layer1 n1_83 (data, 83, layer1_output[83]);
    neuron_layer1 n1_84 (data, 84, layer1_output[84]);
    neuron_layer1 n1_85 (data, 85, layer1_output[85]);
    neuron_layer1 n1_86 (data, 86, layer1_output[86]);
    neuron_layer1 n1_87 (data, 87, layer1_output[87]);
    neuron_layer1 n1_88 (data, 88, layer1_output[88]);
    neuron_layer1 n1_89 (data, 89, layer1_output[89]);
    neuron_layer1 n1_90 (data, 90, layer1_output[90]);
    neuron_layer1 n1_91 (data, 91, layer1_output[91]);
    neuron_layer1 n1_92 (data, 92, layer1_output[92]);
    neuron_layer1 n1_93 (data, 93, layer1_output[93]);
    neuron_layer1 n1_94 (data, 94, layer1_output[94]);
    neuron_layer1 n1_95 (data, 95, layer1_output[95]);
    neuron_layer1 n1_96 (data, 96, layer1_output[96]);
    neuron_layer1 n1_97 (data, 97, layer1_output[97]);
    neuron_layer1 n1_98 (data, 98, layer1_output[98]);
    neuron_layer1 n1_99 (data, 99, layer1_output[99]);
    neuron_layer1 n1_100 (data, 100, layer1_output[100]);
    neuron_layer1 n1_101 (data, 101, layer1_output[101]);
    neuron_layer1 n1_102 (data, 102, layer1_output[102]);
    neuron_layer1 n1_103 (data, 103, layer1_output[103]);
    neuron_layer1 n1_104 (data, 104, layer1_output[104]);
    neuron_layer1 n1_105 (data, 105, layer1_output[105]);
    neuron_layer1 n1_106 (data, 106, layer1_output[106]);
    neuron_layer1 n1_107 (data, 107, layer1_output[107]);
    neuron_layer1 n1_108 (data, 108, layer1_output[108]);
    neuron_layer1 n1_109 (data, 109, layer1_output[109]);
    neuron_layer1 n1_110 (data, 110, layer1_output[110]);
    neuron_layer1 n1_111 (data, 111, layer1_output[111]);
    neuron_layer1 n1_112 (data, 112, layer1_output[112]);
    neuron_layer1 n1_113 (data, 113, layer1_output[113]);
    neuron_layer1 n1_114 (data, 114, layer1_output[114]);
    neuron_layer1 n1_115 (data, 115, layer1_output[115]);
    neuron_layer1 n1_116 (data, 116, layer1_output[116]);
    neuron_layer1 n1_117 (data, 117, layer1_output[117]);
    neuron_layer1 n1_118 (data, 118, layer1_output[118]);
    neuron_layer1 n1_119 (data, 119, layer1_output[119]);
    neuron_layer1 n1_120 (data, 120, layer1_output[120]);
    neuron_layer1 n1_121 (data, 121, layer1_output[121]);
    neuron_layer1 n1_122 (data, 122, layer1_output[122]);
    neuron_layer1 n1_123 (data, 123, layer1_output[123]);
    neuron_layer1 n1_124 (data, 124, layer1_output[124]);
    neuron_layer1 n1_125 (data, 125, layer1_output[125]);
    neuron_layer1 n1_126 (data, 126, layer1_output[126]);
    neuron_layer1 n1_127 (data, 127, layer1_output[127]);
    neuron_layer1 n1_128 (data, 128, layer1_output[128]);
    neuron_layer1 n1_129 (data, 129, layer1_output[129]);
    neuron_layer1 n1_130 (data, 130, layer1_output[130]);
    neuron_layer1 n1_131 (data, 131, layer1_output[131]);
    neuron_layer1 n1_132 (data, 132, layer1_output[132]);
    neuron_layer1 n1_133 (data, 133, layer1_output[133]);
    neuron_layer1 n1_134 (data, 134, layer1_output[134]);
    neuron_layer1 n1_135 (data, 135, layer1_output[135]);
    neuron_layer1 n1_136 (data, 136, layer1_output[136]);
    neuron_layer1 n1_137 (data, 137, layer1_output[137]);
    neuron_layer1 n1_138 (data, 138, layer1_output[138]);
    neuron_layer1 n1_139 (data, 139, layer1_output[139]);
    neuron_layer1 n1_140 (data, 140, layer1_output[140]);
    neuron_layer1 n1_141 (data, 141, layer1_output[141]);
    neuron_layer1 n1_142 (data, 142, layer1_output[142]);
    neuron_layer1 n1_143 (data, 143, layer1_output[143]);
    neuron_layer1 n1_144 (data, 144, layer1_output[144]);
    neuron_layer1 n1_145 (data, 145, layer1_output[145]);
    neuron_layer1 n1_146 (data, 146, layer1_output[146]);
    neuron_layer1 n1_147 (data, 147, layer1_output[147]);
    neuron_layer1 n1_148 (data, 148, layer1_output[148]);
    neuron_layer1 n1_149 (data, 149, layer1_output[149]);
    neuron_layer1 n1_150 (data, 150, layer1_output[150]);
    neuron_layer1 n1_151 (data, 151, layer1_output[151]);
    neuron_layer1 n1_152 (data, 152, layer1_output[152]);
    neuron_layer1 n1_153 (data, 153, layer1_output[153]);
    neuron_layer1 n1_154 (data, 154, layer1_output[154]);
    neuron_layer1 n1_155 (data, 155, layer1_output[155]);
    neuron_layer1 n1_156 (data, 156, layer1_output[156]);
    neuron_layer1 n1_157 (data, 157, layer1_output[157]);
    neuron_layer1 n1_158 (data, 158, layer1_output[158]);
    neuron_layer1 n1_159 (data, 159, layer1_output[159]);
    neuron_layer1 n1_160 (data, 160, layer1_output[160]);
    neuron_layer1 n1_161 (data, 161, layer1_output[161]);
    neuron_layer1 n1_162 (data, 162, layer1_output[162]);
    neuron_layer1 n1_163 (data, 163, layer1_output[163]);
    neuron_layer1 n1_164 (data, 164, layer1_output[164]);
    neuron_layer1 n1_165 (data, 165, layer1_output[165]);
    neuron_layer1 n1_166 (data, 166, layer1_output[166]);
    neuron_layer1 n1_167 (data, 167, layer1_output[167]);
    neuron_layer1 n1_168 (data, 168, layer1_output[168]);
    neuron_layer1 n1_169 (data, 169, layer1_output[169]);
    neuron_layer1 n1_170 (data, 170, layer1_output[170]);
    neuron_layer1 n1_171 (data, 171, layer1_output[171]);
    neuron_layer1 n1_172 (data, 172, layer1_output[172]);
    neuron_layer1 n1_173 (data, 173, layer1_output[173]);
    neuron_layer1 n1_174 (data, 174, layer1_output[174]);
    neuron_layer1 n1_175 (data, 175, layer1_output[175]);
    neuron_layer1 n1_176 (data, 176, layer1_output[176]);
    neuron_layer1 n1_177 (data, 177, layer1_output[177]);
    neuron_layer1 n1_178 (data, 178, layer1_output[178]);
    neuron_layer1 n1_179 (data, 179, layer1_output[179]);
    neuron_layer1 n1_180 (data, 180, layer1_output[180]);
    neuron_layer1 n1_181 (data, 181, layer1_output[181]);
    neuron_layer1 n1_182 (data, 182, layer1_output[182]);
    neuron_layer1 n1_183 (data, 183, layer1_output[183]);
    neuron_layer1 n1_184 (data, 184, layer1_output[184]);
    neuron_layer1 n1_185 (data, 185, layer1_output[185]);
    neuron_layer1 n1_186 (data, 186, layer1_output[186]);
    neuron_layer1 n1_187 (data, 187, layer1_output[187]);
    neuron_layer1 n1_188 (data, 188, layer1_output[188]);
    neuron_layer1 n1_189 (data, 189, layer1_output[189]);
    neuron_layer1 n1_190 (data, 190, layer1_output[190]);
    neuron_layer1 n1_191 (data, 191, layer1_output[191]);
    neuron_layer1 n1_192 (data, 192, layer1_output[192]);
    neuron_layer1 n1_193 (data, 193, layer1_output[193]);
    neuron_layer1 n1_194 (data, 194, layer1_output[194]);
    neuron_layer1 n1_195 (data, 195, layer1_output[195]);
    neuron_layer1 n1_196 (data, 196, layer1_output[196]);
    neuron_layer1 n1_197 (data, 197, layer1_output[197]);
    neuron_layer1 n1_198 (data, 198, layer1_output[198]);
    neuron_layer1 n1_199 (data, 199, layer1_output[199]);

    neuron_layer2 n2_0 (layer1_output, 0, layer2_output[0]);
    neuron_layer2 n2_1 (layer1_output, 1, layer2_output[1]);
    neuron_layer2 n2_2 (layer1_output, 2, layer2_output[2]);
    neuron_layer2 n2_3 (layer1_output, 3, layer2_output[3]);
    neuron_layer2 n2_4 (layer1_output, 4, layer2_output[4]);
    neuron_layer2 n2_5 (layer1_output, 5, layer2_output[5]);
    neuron_layer2 n2_6 (layer1_output, 6, layer2_output[6]);
    neuron_layer2 n2_7 (layer1_output, 7, layer2_output[7]);
    neuron_layer2 n2_8 (layer1_output, 8, layer2_output[8]);
    neuron_layer2 n2_9 (layer1_output, 9, layer2_output[9]);
    neuron_layer2 n2_10 (layer1_output, 10, layer2_output[10]);
    neuron_layer2 n2_11 (layer1_output, 11, layer2_output[11]);
    neuron_layer2 n2_12 (layer1_output, 12, layer2_output[12]);
    neuron_layer2 n2_13 (layer1_output, 13, layer2_output[13]);
    neuron_layer2 n2_14 (layer1_output, 14, layer2_output[14]);
    neuron_layer2 n2_15 (layer1_output, 15, layer2_output[15]);
    neuron_layer2 n2_16 (layer1_output, 16, layer2_output[16]);
    neuron_layer2 n2_17 (layer1_output, 17, layer2_output[17]);
    neuron_layer2 n2_18 (layer1_output, 18, layer2_output[18]);
    neuron_layer2 n2_19 (layer1_output, 19, layer2_output[19]);
    neuron_layer2 n2_20 (layer1_output, 20, layer2_output[20]);
    neuron_layer2 n2_21 (layer1_output, 21, layer2_output[21]);
    neuron_layer2 n2_22 (layer1_output, 22, layer2_output[22]);
    neuron_layer2 n2_23 (layer1_output, 23, layer2_output[23]);
    neuron_layer2 n2_24 (layer1_output, 24, layer2_output[24]);
    neuron_layer2 n2_25 (layer1_output, 25, layer2_output[25]);
    neuron_layer2 n2_26 (layer1_output, 26, layer2_output[26]);
    neuron_layer2 n2_27 (layer1_output, 27, layer2_output[27]);
    neuron_layer2 n2_28 (layer1_output, 28, layer2_output[28]);
    neuron_layer2 n2_29 (layer1_output, 29, layer2_output[29]);
    neuron_layer2 n2_30 (layer1_output, 30, layer2_output[30]);
    neuron_layer2 n2_31 (layer1_output, 31, layer2_output[31]);
    neuron_layer2 n2_32 (layer1_output, 32, layer2_output[32]);
    neuron_layer2 n2_33 (layer1_output, 33, layer2_output[33]);
    neuron_layer2 n2_34 (layer1_output, 34, layer2_output[34]);
    neuron_layer2 n2_35 (layer1_output, 35, layer2_output[35]);
    neuron_layer2 n2_36 (layer1_output, 36, layer2_output[36]);
    neuron_layer2 n2_37 (layer1_output, 37, layer2_output[37]);
    neuron_layer2 n2_38 (layer1_output, 38, layer2_output[38]);
    neuron_layer2 n2_39 (layer1_output, 39, layer2_output[39]);
    neuron_layer2 n2_40 (layer1_output, 40, layer2_output[40]);
    neuron_layer2 n2_41 (layer1_output, 41, layer2_output[41]);
    neuron_layer2 n2_42 (layer1_output, 42, layer2_output[42]);
    neuron_layer2 n2_43 (layer1_output, 43, layer2_output[43]);
    neuron_layer2 n2_44 (layer1_output, 44, layer2_output[44]);
    neuron_layer2 n2_45 (layer1_output, 45, layer2_output[45]);
    neuron_layer2 n2_46 (layer1_output, 46, layer2_output[46]);
    neuron_layer2 n2_47 (layer1_output, 47, layer2_output[47]);
    neuron_layer2 n2_48 (layer1_output, 48, layer2_output[48]);
    neuron_layer2 n2_49 (layer1_output, 49, layer2_output[49]);

    neuron_layer3 n3_0 (layer2_output, 0, result[0]);
    neuron_layer3 n3_1 (layer2_output, 1, result[1]);
    neuron_layer3 n3_2 (layer2_output, 2, result[2]);
    neuron_layer3 n3_3 (layer2_output, 3, result[3]);
    neuron_layer3 n3_4 (layer2_output, 4, result[4]);
    neuron_layer3 n3_5 (layer2_output, 5, result[5]);
    neuron_layer3 n3_6 (layer2_output, 6, result[6]);
    neuron_layer3 n3_7 (layer2_output, 7, result[7]);
    neuron_layer3 n3_8 (layer2_output, 8, result[8]);
    neuron_layer3 n3_9 (layer2_output, 9, result[9]);


endmodule // network

module network (picture);
    input logic [767:0] picture;

endmodule // network

module neuron(input [0:15] bias);
    for(int i = 0; i < )

endmodule // neuron
